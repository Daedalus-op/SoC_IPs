`ifndef UART_SETTINGS
  `define UART_SETTINGS

//  `define DMA_SUPPORT // Enable DMA ports
//  `define PERI8 // 8 bit peripheral, Work in progress 

`endif
